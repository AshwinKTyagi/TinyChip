
module alu (
	input logic bit_type
	input logic[N-1:0] operand1, operand2,
	input logic[3:0] operation,
	output logic[(2*N)-1:0] alu_out
)

	//bit_type

endmodule: alu