module register_file



